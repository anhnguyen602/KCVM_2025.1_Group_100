module test_ALU();

parameter ADD_A_SIZE = 1000;
parameter ADD_B_SIZE = 1000;
parameter ADD_C_SIZE = 1000;
parameter ADD_Cout_SIZE = 1000;
parameter ADD_A_WIDTH = 32;
parameter ADD_B_WIDTH = 32;
parameter ADD_C_WIDTH = 32;
parameter ADD_Cout_WIDTH = 1;

parameter SUB_A_SIZE = 1000;
parameter SUB_B_SIZE = 1000;
parameter SUB_C_SIZE = 1000;
parameter SUB_Cout_SIZE = 1000;
parameter SUB_A_WIDTH = 32;
parameter SUB_B_WIDTH = 32;
parameter SUB_C_WIDTH = 32;
parameter SUB_Cout_WIDTH = 1;

parameter MUL_M_SIZE = 1000;
parameter MUL_Q_SIZE = 1000;
parameter MUL_A_SIZE = 1000;
parameter MUL_M_WIDTH = 32;
parameter MUL_Q_WIDTH = 32;
parameter MUL_A_WIDTH = 64;

parameter DIV_Z_SIZE = 1000;
parameter DIV_D_SIZE = 1000;
parameter DIV_Q_SIZE = 1000;
parameter DIV_R_SIZE = 1000;
parameter DIV_Z_WIDTH = 64;
parameter DIV_D_WIDTH = 32;
parameter DIV_Q_WIDTH = 32;
parameter DIV_R_WIDTH = 32;

parameter INPUT_A_32        = "./input_data/ADD&SUB_input_A.txt";
parameter INPUT_B_32        = "./input_data/ADD&SUB_input_B.txt";
parameter OUTPUT_C_ADD      = "./input_data/ADD_output_C.txt";
parameter OUTPUT_Cout_ADD   = "./input_data/ADD_output_Cout.txt";
parameter OUTPUT_C_SUB      = "./input_data/SUB_output_C.txt";
parameter OUTPUT_Cout_SUB   = "./input_data/SUB_output_Cout.txt";

parameter INPUT_M_MUL       = "./input_data/MUL_input_M.txt";
parameter INPUT_Q_MUL       = "./input_data/MUL_input_Q.txt";
parameter OUTPUT_A_MUL      = "./input_data/MUL_output_A.txt";

parameter INPUT_Z_DIV       = "./input_data/DIV_input_Z.txt";
parameter INPUT_D_DIV       = "./input_data/DIV_input_D.txt";
parameter OUTPUT_Q_DIV      = "./input_data/DIV_output_Q.txt";
parameter OUTPUT_R_DIV      = "./input_data/DIV_output_R.txt";
parameter OUTPUT_FLAG_OVERFLOW_DIV = "./input_data/DIV_flag_overflow.txt";

reg clk;
always #1 clk = ~clk;
initial begin
    clk = 0;
end
reg reset;
reg en;

reg signed [ADD_A_WIDTH-1:0] ADD_input_A [0:(ADD_A_SIZE-1)];
reg signed [ADD_B_WIDTH-1:0] ADD_input_B [0:(ADD_B_SIZE-1)];
reg signed [ADD_C_WIDTH-1:0] ADD_output_C [0:(ADD_C_SIZE-1)];
reg signed ADD_output_Cout [0:(ADD_Cout_SIZE-1)];

reg signed [SUB_A_WIDTH-1:0] SUB_input_A [0:(SUB_A_SIZE-1)];
reg signed [SUB_B_WIDTH-1:0] SUB_input_B [0:(SUB_B_SIZE-1)];
reg signed [SUB_C_WIDTH-1:0] SUB_output_C [0:(SUB_C_SIZE-1)];
reg signed SUB_output_Cout [0:(SUB_Cout_SIZE-1)];

reg signed [MUL_M_WIDTH-1:0] MUL_input_M [0:(MUL_M_SIZE-1)];
reg signed [MUL_Q_WIDTH-1:0] MUL_input_Q [0:(MUL_Q_SIZE-1)];
reg signed [MUL_A_WIDTH-1:0] MUL_output_A [0:(MUL_A_SIZE-1)];

reg signed [DIV_Z_WIDTH-1:0] DIV_input_Z [0:(DIV_Z_SIZE-1)];
reg signed [DIV_D_WIDTH-1:0] DIV_input_D [0:(DIV_D_SIZE-1)];
reg signed [DIV_Q_WIDTH-1:0] DIV_output_Q [0:(DIV_Q_SIZE-1)];
reg signed [DIV_R_WIDTH-1:0] DIV_output_R [0:(DIV_R_SIZE-1)];
reg DIV_flag_overflow [0:(DIV_R_SIZE-1)];

// reg signed [ADD_A_WIDTH-1:0] ADD_DUT_input_A;
// reg signed [ADD_B_WIDTH-1:0] ADD_DUT_input_B;
// wire signed [ADD_C_WIDTH-1:0] ADD_DUT_output_C;
// wire signed ADD_DUT_output_Cout;

// reg signed [SUB_A_WIDTH-1:0] SUB_DUT_input_A;
// reg signed [SUB_B_WIDTH-1:0] SUB_DUT_input_B;
// wire signed [SUB_C_WIDTH-1:0] SUB_DUT_output_C;
// wire signed SUB_DUT_output_Cout;

reg signed [MUL_M_WIDTH-1:0] MUL_DUT_input_M;
reg signed [MUL_Q_WIDTH-1:0] MUL_DUT_input_Q;
wire signed [MUL_A_WIDTH-1:0] MUL_DUT_output_A;
wire MUL_DUT_done;

// reg signed [DIV_Z_WIDTH-1:0] DIV_DUT_input_Z;
// reg signed [DIV_D_WIDTH-1:0] DIV_DUT_input_D;
// wire signed [DIV_Q_WIDTH-1:0] DIV_DUT_output_Q;
// wire signed [DIV_R_WIDTH-1:0] DIV_DUT_output_R;
// wire DIV_DUT_done;
// wire [3:0] DIV_DUT_flag;
// parameter OVERFLOW_BIT = 3;

reg signed [31:0] ALU_DUT_num_1;
reg signed [31:0] ALU_DUT_num_2;
reg signed [31:0] ALU_DUT_sub_reg_input;
reg signed [3:0] ALU_DUT_opcode;
wire signed [31:0] ALU_DUT_result;
wire signed [31:0] ALU_DUT_sub_reg_result;
wire signed ALU_DUT_done;
wire signed [3:0] ALU_DUT_flag;
wire  signed  [63:0] ALU_DUT_MUL_result = {ALU_DUT_sub_reg_result, ALU_DUT_result};
reg   signed [63:0] ALU_DUT_DIV_Z;
wire  signed  [31:0] ALU_DUT_DIV_sub_reg_input = ALU_DUT_DIV_Z[63:32];
wire  signed  [31:0] ALU_DUT_DIV_num_1 = ALU_DUT_DIV_Z[31:0];

    ALU #(.WIDTH(32)) ALU_DUT(
        .num_1(ALU_DUT_num_1),
        .num_2(ALU_DUT_num_2),
        .sub_reg_input(ALU_DUT_sub_reg_input),
        .opcode(ALU_DUT_opcode),
        .result(ALU_DUT_result),
        .sub_reg_result(ALU_DUT_sub_reg_result),
        .clk(clk),
        .flag(ALU_DUT_flag),
        .done(ALU_DUT_done)
    );

    integer i;
    integer ADD_ERROR = 0;
    integer SUB_ERROR = 0;
    integer NEG_ERROR = 0;
    integer MUL_ERROR = 0;
    integer DIV_ERROR = 0;
    integer AND_ERROR = 0;
    integer OR_ERROR = 0;
    integer XOR_ERROR = 0;
    integer NOT_ERROR = 0;

    parameter ADD = 4'b0000;
    parameter SUB = 4'b0001;
    parameter MUL = 4'b0010;
    parameter DIV = 4'b0011; // chú ý trường hợp chia cho 0
    parameter NEG = 4'b0100; // bù 2 của num_1
    parameter AND = 4'b0101;
    parameter OR  = 4'b0110;
    parameter XOR = 4'b0111;
    parameter NOT = 4'b1000; // đảo của num_1

    parameter OVERFLOW=3;
    parameter ZERO=2;
    parameter SIGN=1;
    parameter CARRY=0;


// /* // ALU TEST_____________________________________________________________________________________________________
initial begin
    clk = 0;
    reset = 1;
    en = 0;
// 
    $readmemh(INPUT_A_32, ADD_input_A);
    $readmemh(INPUT_B_32, ADD_input_B);
    $readmemh(OUTPUT_C_ADD, ADD_output_C);
    $readmemh(OUTPUT_Cout_ADD, ADD_output_Cout);

    $readmemh(INPUT_A_32, SUB_input_A);
    $readmemh(INPUT_B_32, SUB_input_B);
    $readmemh(OUTPUT_C_SUB, SUB_output_C);
    $readmemh(OUTPUT_Cout_SUB, SUB_output_Cout);

    $readmemh(INPUT_M_MUL, MUL_input_M);
    $readmemh(INPUT_Q_MUL, MUL_input_Q);
    $readmemh(OUTPUT_A_MUL, MUL_output_A);

    $readmemh(INPUT_Z_DIV, DIV_input_Z);
    $readmemh(INPUT_D_DIV, DIV_input_D);
    $readmemh(OUTPUT_Q_DIV, DIV_output_Q);
    $readmemh(OUTPUT_R_DIV, DIV_output_R);
    $readmemh(OUTPUT_FLAG_OVERFLOW_DIV, DIV_flag_overflow);
// 
// /*

    ALU_DUT_opcode = ADD;

    for(i = 0; i < ADD_A_SIZE; i = i + 1) begin
        #1;
            ALU_DUT_num_1 = ADD_input_A[i];
            ALU_DUT_num_2 = ADD_input_B[i];
        #3;
        while(ALU_DUT_done == 0) begin
            #1;
        end
        if(ALU_DUT_result != ADD_output_C[i] || ALU_DUT_flag[CARRY] != ADD_output_Cout[i]) begin
            if(ALU_DUT_result != ADD_output_Cout[i]) begin
                ADD_ERROR = ADD_ERROR + 1;
                // $display("%t ADD test failed at %d line",$time, i+1);
                // $display("Input: %d + %d = %d Carry out %b", ALU_DUT_num_1, ALU_DUT_num_2, ALU_DUT_result, ALU_DUT_flag[CARRY]);
                // $display("Expected output: %d %d", ADD_output_C[i], ADD_output_Cout[i]);
            end else if (ALU_DUT_flag[CARRY] == 0) begin // không bị overflow
                ADD_ERROR = ADD_ERROR + 1;
                // $display("%t ADD test failed at %d line (NO Carry out)",$time, i+1);
                // $display("Input: %h + %h = %h Carry out %b", ADD_DUT_input_A, ADD_DUT_input_B, ADD_DUT_output_C, ADD_DUT_output_Cout);
                // $display("Expected output: %h %h", ADD_output_C[i], ADD_output_Cout[i]);
            end
        end
        #2;
    end
    if(ADD_ERROR == 0) begin
        $display("______________________________________________ADD test passed___________________________________________");
    end else begin
        $display("___________________________________________ADD passed %d/%d test cases___________________________________", ADD_A_SIZE - ADD_ERROR, ADD_A_SIZE);
    end
// * /

    ALU_DUT_opcode = SUB;

    for(i = 0; i < SUB_A_SIZE; i = i + 1) begin
        #1;
            ALU_DUT_num_1 = SUB_input_A[i];
            ALU_DUT_num_2 = SUB_input_B[i];
        #3;
        while(ALU_DUT_done == 0) begin
            #1;
        end
        if(ALU_DUT_result != SUB_output_C[i] || ALU_DUT_flag[CARRY] != SUB_output_Cout[i]) begin
            if(ALU_DUT_result != SUB_output_Cout[i]) begin
                SUB_ERROR = SUB_ERROR + 1;
                // $display("%t SUB test failed at %d line",$time, i+1);
                // $display("Input: %d + %d = %d Carry out %b", ALU_DUT_num_1, ALU_DUT_num_2, ALU_DUT_result, ALU_DUT_flag[CARRY]);
                // $display("Expected output: %d %d", SUB_output_C[i], SUB_output_Cout[i]);
            end else if (ALU_DUT_flag[CARRY] == 0) begin // không bị overflow
                SUB_ERROR = SUB_ERROR + 1;
                // $display("%t SUB test failed at %d line (NO Carry out)",$time, i+1);
                // $display("Input: %h + %h = %h Carry out %b", SUB_DUT_input_A, SUB_DUT_input_B, SUB_DUT_output_C, SUB_DUT_output_Cout);
                // $display("Expected output: %h %h", SUB_output_C[i], ADD_output_Cout[i]);
            end
        end
        #2;
    end

    if(SUB_ERROR == 0) begin
        $display("______________________________________________SUB test passed___________________________________________");
    end else begin
        $display("___________________________________________SUB passed %d/%d test cases___________________________________", SUB_A_SIZE - SUB_ERROR, SUB_A_SIZE);
    end

//
// /*
    #3;
    ALU_DUT_opcode = MUL;

    for(i = 0; i < MUL_M_SIZE; i = i + 1) begin
        ALU_DUT_num_1 = MUL_input_M[i];
        ALU_DUT_num_2 = MUL_input_Q[i];
        #2;
        while(ALU_DUT_done == 0) begin
            #1;
        end
        #1;
        if(ALU_DUT_MUL_result != MUL_output_A[i]) begin
            MUL_ERROR = MUL_ERROR + 1;
            // $display("%t MUL test failed at %d line",$time, i+1);
            // $display("Input: %b * %b = %b", ALU_DUT_num_1, ALU_DUT_num_2, ALU_DUT_MUL_result);
            // $display("Expected output: %b", MUL_output_A[i]);
        end
    end

    if(MUL_ERROR == 0) begin
        $display("______________________________________________MUL test passed___________________________________________");
    end else begin
        $display("___________________________________________MUL passed %d/%d test cases___________________________________", MUL_M_SIZE - MUL_ERROR, MUL_M_SIZE);
    end
// / //
    #4;

    ALU_DUT_opcode = DIV;

    // /*
    // DIV_DUT_input_Z = DIV_input_Z[0];
    // DIV_DUT_input_D = DIV_input_D[0];
            // $display("DIV_DUT_input_Z = %h, DIV_DUT_input_D = %h, INPUT DATA: %h %h\n", DIV_DUT_input_Z, DIV_DUT_input_D, DIV_input_Z[0], DIV_input_D[0]);
    i = 0;
    for(i = 0; i < DIV_Z_SIZE; i = i + 1) begin
        // if(ALU_DUT_done == 1) begin

            ALU_DUT_DIV_Z = DIV_input_Z[i]; 
            #1;
            ALU_DUT_sub_reg_input = ALU_DUT_DIV_sub_reg_input;
            ALU_DUT_num_1 = ALU_DUT_DIV_num_1;
            ALU_DUT_num_2 = DIV_input_D[i];      
        // end
        #2;
            // $display("DIV_DUT_input_Z = %h, DIV_DUT_input_D = %h, INPUT DATA: %h %h\n", DIV_DUT_input_Z, DIV_DUT_input_D, DIV_input_Z[i], DIV_input_D[i]);
            // #1;
        while(ALU_DUT_done == 0) begin
            // $display (" %t i = %d DIV_DUT_done = %d CALCULATING...",$time, i, DIV_DUT_done);
            // $display("CALCULATING...");
            #1;
        end

        if(ALU_DUT_result != DIV_output_Q[i] || ALU_DUT_sub_reg_result != DIV_output_R[i] || ALU_DUT_flag[OVERFLOW] != DIV_flag_overflow[i])   begin
            if(ALU_DUT_flag[OVERFLOW] != DIV_flag_overflow[i]) begin
                DIV_ERROR = DIV_ERROR + 1;
                // $display("%t DIV test failed at i = %d, at %d line, Expected OVERFLOW = %d",$time, i, i+1, DIV_flag_overflow[i]);
                // $display("DUT output: %h (%d) / %h (%d) = %h (%d) R %h (%d), OVERFLOW = %d", ALU_DUT_DIV_Z, ALU_DUT_DIV_Z, ALU_DUT_num_2, ALU_DUT_num_2, ALU_DUT_result, ALU_DUT_result, ALU_DUT_sub_reg_result, ALU_DUT_sub_reg_result, ALU_DUT_flag[OVERFLOW]);
                // $display("Expected output: Q =  %h (%d); R = %h (%d), OVERFLOW = %d", DIV_output_Q[i], DIV_output_Q[i], DIV_output_R[i], DIV_output_R[i], DIV_flag_overflow[i]);
            end else if(DIV_flag_overflow[i] == 0) begin
                DIV_ERROR = DIV_ERROR + 1;
                // $display("%t DIV test failed at i = %d, at %d line (NO OVERFLOW)",$time, i, i+1);
                // $display("DUT output: %h (%d) / %h (%d) = %h (%d) R %h (%d), OVERFLOW = %d", ALU_DUT_DIV_Z, ALU_DUT_DIV_Z, ALU_DUT_num_2, ALU_DUT_num_2, ALU_DUT_result, ALU_DUT_result, ALU_DUT_sub_reg_result, ALU_DUT_sub_reg_result, ALU_DUT_flag[OVERFLOW]);
                // $display("Expected output: Q =  %h (%d); R = %h (%d), OVERFLOW = %d", DIV_output_Q[i], DIV_output_Q[i], DIV_output_R[i], DIV_output_R[i], DIV_flag_overflow[i]);
            end
        end
    end

    if(DIV_ERROR == 0) begin
        $display("______________________________________________DIV test passed___________________________________________");
    end else begin
        $display("___________________________________________DIV passed %d/%d test cases___________________________________", DIV_Z_SIZE - DIV_ERROR, DIV_Z_SIZE);
    end
//
    $finish;

end
// */

// reg en;

// mul MUL_DUT(
//     .M_in(MUL_DUT_input_M),
//     .Q_in(MUL_DUT_input_Q),
//     .clk(clk),
//     .reset(reset),
//     .en(en),
//     .done(MUL_DUT_done),
//     .A_out(MUL_DUT_output_A)
// );


// initial begin
//     clk = 0;
//     reset = 1;
//     en = 0;
// // 
//     $readmemh(INPUT_A_32, ADD_input_A);
//     $readmemh(INPUT_B_32, ADD_input_B);
//     $readmemh(OUTPUT_C_ADD, ADD_output_C);
//     $readmemh(OUTPUT_Cout_ADD, ADD_output_Cout);

//     $readmemh(INPUT_A_32, SUB_input_A);
//     $readmemh(INPUT_B_32, SUB_input_B);
//     $readmemh(OUTPUT_C_SUB, SUB_output_C);
//     $readmemh(OUTPUT_Cout_SUB, SUB_output_Cout);

//     $readmemh(INPUT_M_MUL, MUL_input_M);
//     $readmemh(INPUT_Q_MUL, MUL_input_Q);
//     $readmemh(OUTPUT_A_MUL, MUL_output_A);

//     $readmemh(INPUT_Z_DIV, DIV_input_Z);
//     $readmemh(INPUT_D_DIV, DIV_input_D);
//     $readmemh(OUTPUT_Q_DIV, DIV_output_Q);
//     $readmemh(OUTPUT_R_DIV, DIV_output_R);
//     $readmemh(OUTPUT_FLAG_OVERFLOW_DIV, DIV_flag_overflow);
// //  
//     #3;
//     reset = 0;
//     en = 1;
//     for(i = 0; i < MUL_M_SIZE; i = i + 1) begin
//         MUL_DUT_input_M = MUL_input_M[i];
//         MUL_DUT_input_Q = MUL_input_Q[i];
//         #1;
//         while(MUL_DUT_done == 0) begin
//             #1;
//         end
//         #1;
//         if(MUL_DUT_output_A != MUL_output_A[i]) begin
//             MUL_ERROR = MUL_ERROR + 1;
//             $display("%t MUL test failed at %d line",$time, i+1);
//             $display("Input: %b (%d) * %b (%d) = %b (%d)", MUL_DUT_input_M, MUL_DUT_input_M, MUL_DUT_input_Q, MUL_DUT_input_Q,  MUL_DUT_output_A, MUL_DUT_output_A);
//             $display("Expected output: %b (%d)", MUL_output_A[i], MUL_output_A[i]);
//             $display("%b", (MUL_output_A[i] ^ MUL_DUT_output_A));
//         end else begin
//             // $display("%t MUL test passed at %d line",$time, i+1);
//             // $display("Input: %h * %h = %h", MUL_DUT_input_M, MUL_DUT_input_Q, MUL_DUT_output_A);
//         end
//     end

//     if(MUL_ERROR == 0) begin
//         $display("______________________________________________MUL test passed___________________________________________");
//     end else begin
//         $display("___________________________________________MUL passed %d/%d test cases___________________________________", MUL_M_SIZE - MUL_ERROR, MUL_M_SIZE);
//     end

//     $finish;

// end


    always @(ALU_DUT_MUL_result, ALU_DUT_flag) begin
        if(ALU_DUT_opcode == MUL && ALU_DUT_done)
        $display("Num 1 = %d, num 2 = %d, result = %d, flag = %b", ALU_DUT_num_1, ALU_DUT_num_2, ALU_DUT_MUL_result, ALU_DUT_flag);
    end

endmodule


// 10000000000000000000000000000000 * 10010011011001010101100110111010 = 0011011001001101010100110010000100000000000000000000000000000000

// 10000000000000000000000000000000 (-2147483648) * 10010011011001010101100110111010 (-1822074438)

// 0011011001001101010100110010001100000000000000000000000000000000 (  3912875061043789824)
// 0011011001001101010100110010000100000000000000000000000000000000

/*
# 0000000000000000000000000000111100000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000011111100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000001111000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000011111100000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000111100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000111100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000111100000000000000000000000000000000
# 0000000000000000000000000000011100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000001111000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000111000000000000000000000000000000000
# 0000000000000000000000000000111100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000001111100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000011100000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000011111000000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000001111111000000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000111111100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000011100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000111100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000111100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000001111000000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000011100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000011100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000011100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000011100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000111100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000111100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000011100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000011100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000111000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000011100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000011100000000000000000000000000000000
# 0000000000000000000000001111111100000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000011111111000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000011100000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000111100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000111000000000000000000000000000000000
# 0000000000000000000000000001111100000000000000000000000000000000
# 0000000000000000000000000000111000000000000000000000000000000000
# 0000000000000000000000000000111100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000011100000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000
# 0000000000000000000000000000011100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000000100000000000000000000000000000000
# 0000000000000000000000000000001100000000000000000000000000000000
# 0000000000000000000000000000011000000000000000000000000000000000
# 0000000000000000000000000000001000000000000000000000000000000000

10000000000000000000000000000000 (-2147483648) * 100 010 001 110 011 100 011 011 011 011 100 011 101 111 101 100 (-1822074438)

100     010     001     110     011     100     010     010     010     011     100     011     101     111     101     100

-2M     M      M        -M      2M     -2M      M       M        M      2M       -2M     2M     -M       0       -M     -2M

// */